module name(
    port_list
);
    begin
        if(cong) {
            stop
        }
    end
endmodule